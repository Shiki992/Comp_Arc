`include "c432.v"
module ctest();
reg N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
wire N223,N329,N370,N421,N430,N431,N432;
c432 HA01(N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,
	initial
		begin
N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,=0;
#5 N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,=0;	
end
initial
		$monitor($time,"N1,n4,n8,n11,n14,n17,n21,n24,n27,n30,=%b N223,n329,n370,n421,n430,n431,n432;=%b ",N1,N4,N8,N11,N14,N17,N21,N24,N27,N30,,N223,N329,N370,N421,N430,N431,N432;,);
endmodule