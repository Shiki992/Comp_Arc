`include "fpad.v";
module top();


endmodule /op
