`include "16BA.v"
module sixteentest;
