`include "c17.v"
module ctest();
reg N1,N2,N3,N6,N7;
wire N22,N23;
c17 HA01(N1,N2,N3,N6,N7,N22,N23);
	initial
		begin
N1=0;
N2=0;
N3=0;
N6=0;
N7=0;
#5 N1=0;	N2=1;	N3=0;	N6=1;	N7=1;	
#5 N1=0;	N2=0;	N3=0;	N6=1;	N7=1;	
#5 N1=0;	N2=0;	N3=1;	N6=1;	N7=0;	
#5 N1=0;	N2=0;	N3=1;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
#5 N1=0;	N2=0;	N3=0;	N6=0;	N7=0;	
end
initial
		$monitor($time,"N1=%b N2=%b N3=%b N6=%b N7=%b N22=%b N23=%b ",N1,N2,N3,N6,N7,N22,N23,);
endmodule